module clockctlr(clk_in, clk_out);

input clk_in;
output wire clk_out;

assign clk_out = clk_in;

endmodule
