130101FD 23268102 13040103 232604FE 
232404FE 232204FE 232004FE 232E04FC 
232C04FC 232A04FC 8327C4FE 93871700 
2326F4FE 0327C4FE 9307C003 B377F702 
2324F4FE 0327C4FE 9307C003 B357F702 
13870700 9307C003 B367F702 2322F4FE 
0327C4FE B7170000 938707E1 B357F702 
13870700 93078001 B367F702 2320F4FE 
0327C4FE B7570100 93870718 B357F702 
13870700 9307F001 B367F702 232EF4FC 
0327C4FE B7E72800 938707E8 B357F702 
13870700 9307C000 B367F702 232CF4FC 
0327C4FE B777EA01 938707E0 B357F702 
232AF4FC 6FF05FF5 
